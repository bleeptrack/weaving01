# LEF file generated for my_logo
VERSION 5.8 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO my_logo
   CLASS BLOCK ;
   FOREIGN my_logo 0 0 ;
   SIZE 80.000 BY 80.000 ;
   SYMMETRY X Y ;
   SITE unithd ;
   PIN VDD
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT
         LAYER met1 ;
         RECT 0.000 78.000 80.000 80.000 ;
      END
   END VDD
   PIN VSS
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT
         LAYER met1 ;
         RECT 0.000 0.000 80.000 2.000 ;
      END
   END VSS
   PIN in1
      DIRECTION INPUT ;
      USE SIGNAL ;
      PORT
         LAYER met1 ;
         RECT 2.000 2.000 3.000 3.000 ;
      END
   END in1
   PIN out1
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      PORT
         LAYER met1 ;
         RECT 77.000 77.000 78.000 78.000 ;
      END
   END out1
   OBS
      LAYER met1 ;
      RECT 0.000 0.000 80.000 80.000 ;
   END
END my_logo
