# LEF file generated for FIRST
VERSION 5.8 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

LAYER metal1
   TYPE ROUTING ;
   WIDTH 0.1 ;
   SPACING 0.1 ;
END metal1

LAYER metal2
   TYPE ROUTING ;
   WIDTH 0.1 ;
   SPACING 0.1 ;
END metal2

MACRO FIRST
   CLASS CORE ;
   FOREIGN FIRST 0 0 ;
   SIZE 80.000 BY 80.000 ;
   SYMMETRY X Y ;
   PIN VDD
      DIRECTION INOUT ;
      USE POWER ;
      PORT
         LAYER metal1 ;
         RECT 0.000 79.000 1.000 80.000 ;
      END
   END VDD
   PIN VSS
      DIRECTION INOUT ;
      USE GROUND ;
      PORT
         LAYER metal1 ;
         RECT 0.000 0.000 1.000 1.000 ;
      END
   END VSS
   PIN in1
      DIRECTION INPUT ;
      USE SIGNAL ;
      PORT
         LAYER metal1 ;
         RECT 2.000 2.000 3.000 3.000 ;
      END
   END in1
   PIN out1
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      PORT
         LAYER metal1 ;
         RECT 77.000 77.000 78.000 78.000 ;
      END
   END out1
   OBS
      LAYER metal1 ;
      RECT 0.000 0.000 80.000 80.000 ;
   END
END FIRST
