# LEF file generated for my_logo
VERSION 5.8 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO my_logo
   CLASS BLOCK ;
   FOREIGN my_logo 0 0 ;
   SIZE 32.000 BY 32.000 ;
   SYMMETRY X Y ;
   PIN dummy
      DIRECTION INOUT ;
      USE SIGNAL ;
      PORT
         LAYER Metal1 ;
         RECT 0.000 0.000 1.000 1.000 ;
      END
   END dummy
END my_logo
