# LEF file generated for FIRST
VERSION 5.8 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO FIRST
   CLASS BLOCK ;
   FOREIGN FIRST 0 0 ;
   SIZE 80.000 BY 80.000 ;
   SYMMETRY X Y ;
   SITE core ;
   PIN VDD
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT
         LAYER metal1 ;
         RECT 0.000 78.000 80.000 80.000 ;
      END
   END VDD
   PIN VSS
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT
         LAYER metal1 ;
         RECT 0.000 0.000 80.000 2.000 ;
      END
   END VSS
   PIN in1
      DIRECTION INPUT ;
      USE SIGNAL ;
      PORT
         LAYER metal1 ;
         RECT 2.000 2.000 3.000 3.000 ;
      END
   END in1
   PIN out1
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      PORT
         LAYER metal1 ;
         RECT 77.000 77.000 78.000 78.000 ;
      END
   END out1
   OBS
      LAYER metal1 ;
      RECT 0.000 0.000 80.000 80.000 ;
   END
END FIRST
