  X �     2�     2 library  >A�7KƧ�9D�/��ZT �     2�     2 
FIRST         ,      �      �  @  �  @  �      �          ,  (m      (m  @  5S  @  5S      (m              ,  E�      E�  @  V�  @  V�      E�              ,  c�      c�  @  v�  @  v�      c�              ,  �      �  @  �>  @  �>      �              ,  �c      �c  @  �]  @  �]      �c              ,  ��  �  ��  �  ��  �  ��  �  ��  �          ,  �x      �x  @  �H  @  �H      �x              , C     C  @ 
�  @ 
�     C              , @  � @  � 8�  � 8�  � @  �          ,  �  @  �  >�  �  >�  �  @  �  @          ,  @  %�  @  7�  >�  7�  >�  %�  @  %�          ,  >�  %�  >�  7�  ]�  7�  ]�  %�  >�  %�          ,  c�  @  c�  >�  v�  >�  v�  @  c�  @          ,  �  @  �  >�  �>  >�  �>  @  �  @          ,  �c  @  �c  >�  �]  >�  �]  @  �c  @          ,  ��  %�  ��  7�  ��  7�  ��  %�  ��  %�          ,  ��  %�  ��  7�  �   7�  �   %�  ��  %�          , C  @ C  >� 
�  >� 
�  @ C  @          , (3  @ (3  >� )�  >� )�  @ (3  @          ,      E%      W  @  W  @  E%      E%          ,  (m  >�  (m  ]�  5S  ]�  5S  >�  (m  >�          ,  >�  E%  >�  W  ]�  W  ]�  E%  >�  E%          ,  c�  >�  c�  ]�  v�  ]�  v�  >�  c�  >�          ,  }   E%  }   W  �@  W  �@  E%  }   E%          ,  �c  >�  �c  ]�  �]  ]�  �]  >�  �c  >�          ,  ĭ  >�  ĭ  ]�  ѓ  ]�  ѓ  >�  ĭ  >�          ,  ��  E%  ��  W  �   W  �   E%  ��  E%          , C  >� C  ]� 
�  ]� 
�  >� C  >�          , (3  >� (3  ]� )�  ]� )�  >� (3  >�          ,  �  ]�  �  }   �  }   �  ]�  �  ]�          ,  (m  ]�  (m  }   5S  }   5S  ]�  (m  ]�          ,  >�  ix  >�  qH  ]�  qH  ]�  ix  >�  ix          ,  ]�  ix  ]�  qH  }   qH  }   ix  ]�  ix          ,  }   ix  }   qH  �@  qH  �@  ix  }   ix          ,  �@  ix  �@  qH  ��  qH  ��  ix  �@  ix          ,  ĭ  ]�  ĭ  }   ѓ  }   ѓ  ]�  ĭ  ]�          ,  �x  ]�  �x  }   �H  }   �H  ]�  �x  ]�          ,  �   ix  �   qH @  qH @  ix  �   ix          , (3  ]� (3  }  )�  }  )�  ]� (3  ]�          ,  �  }   �  �@  �  �@  �  }   �  }           ,  (m  }   (m  �@  5S  �@  5S  }   (m  }           ,  >�  �u  >�  ��  ]�  ��  ]�  �u  >�  �u          ,  c�  }   c�  �@  v�  �@  v�  }   c�  }           ,  �  }   �  �@  �>  �@  �>  }   �  }           ,  �@  �u  �@  ��  ��  ��  ��  �u  �@  �u          ,  ĭ  }   ĭ  �@  ѓ  �@  ѓ  }   ĭ  }           ,  �x  }   �x  �@  �H  �@  �H  }   �x  }           ,  �   �u  �   �� @  �� @  �u  �   �u          , @  �u @  �� 8�  �� 8�  �u @  �u          ,      ��      �  @  �  @  ��      ��          ,  (m  �@  (m  ��  5S  ��  5S  �@  (m  �@          ,  E�  �@  E�  ��  V�  ��  V�  �@  E�  �@          ,  ]�  ��  ]�  �  }   �  }   ��  ]�  ��          ,  }   ��  }   �  �@  �  �@  ��  }   ��          ,  �c  �@  �c  ��  �]  ��  �]  �@  �c  �@          ,  ĭ  �@  ĭ  ��  ѓ  ��  ѓ  �@  ĭ  �@          ,  ��  ��  ��  �  �   �  �   ��  ��  ��          , C  �@ C  �� 
�  �� 
�  �@ C  �@          , (3  �@ (3  �� )�  �� )�  �@ (3  �@          ,  �  ��  �  ��  �  ��  �  ��  �  ��          ,  (m  ��  (m  ��  5S  ��  5S  ��  (m  ��          ,  >�  �8  >�  �  ]�  �  ]�  �8  >�  �8          ,  c�  ��  c�  ��  v�  ��  v�  ��  c�  ��          ,  �  ��  �  ��  �>  ��  �>  ��  �  ��          ,  �c  ��  �c  ��  �]  ��  �]  ��  �c  ��          ,  ��  �8  ��  �  ��  �  ��  �8  ��  �8          ,  ��  �8  ��  �  �   �  �   �8  ��  �8          ,  �   �8  �   � @  � @  �8  �   �8          , (3  �� (3  �� )�  �� )�  �� (3  ��          ,      �e      �[  @  �[  @  �e      �e          ,  (m  ��  (m  �   5S  �   5S  ��  (m  ��          ,  >�  �e  >�  �[  ]�  �[  ]�  �e  >�  �e          ,  c�  ��  c�  �   v�  �   v�  ��  c�  ��          ,  }   �e  }   �[  �@  �[  �@  �e  }   �e          ,  �c  ��  �c  �   �]  �   �]  ��  �c  ��          ,  ĭ  ��  ĭ  �   ѓ  �   ѓ  ��  ĭ  ��          ,  �x  ��  �x  �   �H  �   �H  ��  �x  ��          , C  �� C  �  
�  �  
�  �� C  ��          , (3  �� (3  �  )�  �  )�  �� (3  ��          ,  �  �   � @  � @  �  �   �  �           ,  @  �  @ �  >� �  >�  �  @  �          ,  >�  �  >� �  ]� �  ]�  �  >�  �          ,  ]�  �  ]� �  }  �  }   �  ]�  �          ,  }   �  }  �  �@ �  �@  �  }   �          ,  �@  �  �@ �  �� �  ��  �  �@  �          ,  ĭ  �   ĭ @  ѓ @  ѓ  �   ĭ  �           ,  �x  �   �x @  �H @  �H  �   �x  �           ,  �   �  �  � @ � @  �  �   �          , (3  �  (3 @ )� @ )�  �  (3  �           ,  � @  � 8�  � 8�  � @  � @          ,  @ $�  @ ,�  >� ,�  >� $�  @ $�          ,  >� $�  >� ,�  ]� ,�  ]� $�  >� $�          ,  ]� $�  ]� ,�  }  ,�  }  $�  ]� $�          ,  � @  � 8�  �> 8�  �> @  � @          ,  �c @  �c 8�  �] 8�  �] @  �c @          ,  �� $�  �� ,�  �� ,�  �� $�  �� $�          ,  �x @  �x 8�  �H 8�  �H @  �x @          ,  �  $�  �  ,� @ ,� @ $�  �  $�          , (3 @ (3 8� )� 8� )� @ (3 @           ,  �@  ��  �@  �  ��  �  ��  ��  �@  ��           ,  �c  ��  �c  ��  �]  ��  �]  ��  �c  ��           ,  �c  �@  �c  �#  �]  �#  �]  �@  �c  �@           ,  ��  ��  ��  �  ��  �  ��  ��  ��  ��           ,  ĭ  ��  ĭ  ��  ѓ  ��  ѓ  ��  ĭ  ��           ,  ĭ  �@  ĭ  �#  ѓ  �#  ѓ  �@  ĭ  �@           ,  �x  �@  �x  ��  �H  ��  �H  �@  �x  �@           ,  ��  ��  ��  �  �  �  �  ��  ��  ��           ,  �0  ��  �0  �  �   �  �   ��  �0  ��           ,  �   ��  �   � @  � @  ��  �   ��           , C  �� C  �� 
�  �� 
�  �� C  ��           , C  �@ C  �# 
�  �# 
�  �@ C  �@           , @  �� @  � 8�  � 8�  �� @  ��           , (3  �� (3  �� )�  �� )�  �� (3  ��           , (3  �@ (3  �# )�  �# )�  �@ (3  �@           ,  �@  �8  �@  �  ��  �  ��  �8  �@  �8           ,  �c  ��  �c  ��  �]  ��  �]  ��  �c  ��           ,  �c  ��  �c  �P  �]  �P  �]  ��  �c  ��           ,  ĭ  ��  ĭ  ��  ѓ  ��  ѓ  ��  ĭ  ��           ,  ��  �8  ��  �  ��  �  ��  �8  ��  �8           ,  �{  �8  �{  �  ��  �  ��  �8  �{  �8           ,  �x  ��  �x  ��  �H  ��  �H  ��  �x  ��           ,  ��  �8  ��  �  �  �  �  �8  ��  �8           ,  �0  �8  �0  �  �   �  �   �8  �0  �8           , C  �� C  �� 
�  �� 
�  �� C  ��           ,  �   �8  �   � [  � [  �8  �   �8           , �  �8 �  � @  � @  �8 �  �8           , @  �8 @  � 8�  � 8�  �8 @  �8           , (3  �� (3  �� )�  �� )�  �� (3  ��           , (3  �� (3  �P )�  �P )�  �� (3  ��           ,  �@  �e  �@  �[  ��  �[  ��  �e  �@  �e           ,  �c  �C  �c  �   �]  �   �]  �C  �c  �C           ,  �c  ��  �c  �}  �]  �}  �]  ��  �c  ��           ,  ��  �e  ��  �[  ��  �[  ��  �e  ��  �e           ,  ĭ  �C  ĭ  �   ѓ  �   ѓ  �C  ĭ  �C           ,  ĭ  ��  ĭ  �}  ѓ  �}  ѓ  ��  ĭ  ��           ,  ��  �e  ��  �[  �   �[  �   �e  ��  �e           ,  �x  �C  �x  �   �H  �   �H  �C  �x  �C           ,  �x  ��  �x  �}  �H  �}  �H  ��  �x  ��           ,  �   �e  �   �[ @  �[ @  �e  �   �e           , C  �C C  �  
�  �  
�  �C C  �C           , C  �� C  �} 
�  �} 
�  �� C  ��           , @  �e @  �[ 8�  �[ 8�  �e @  �e           , (3  �C (3  �  )�  �  )�  �C (3  �C           , (3  �� (3  �} )�  �} )�  �� (3  ��           ,  �c  �   �c @  �] @  �]  �   �c  �            ,  �@  �  �@ �  �{ �  �{  �  �@  �           ,  �E  �  �E �  �� �  ��  �  �E  �           ,  ��  �  �� �  �� �  ��  �  ��  �           ,  ĭ �  ĭ @  ѓ @  ѓ �  ĭ �           ,  ĭ  �   ĭ  ��  ѓ  ��  ѓ  �   ĭ  �            ,  ��  �  �� �  �  �  �   �  ��  �           ,  �x �  �x @  �H @  �H �  �x �           ,  �x  �   �x  ��  �H  ��  �H  �   �x  �            , C  �  C @ 
� @ 
�  �  C  �            ,  �   �  �  � [ � [  �  �   �           , �  � � � @ � @  � �  �           , @  � @ � 8� � 8�  � @  �           , (3 � (3 @ )� @ )� � (3 �           , (3  �  (3  �� )�  �� )�  �  (3  �            ,  �@ $�  �@ ,�  �� ,�  �� $�  �@ $�           ,  �c 0�  �c 8�  �] 8�  �] 0�  �c 0�           ,  �c @  �c !  �] !  �] @  �c @           ,  ĭ @  ĭ 8�  ѓ 8�  ѓ @  ĭ @           ,  �� $�  �� ,�  �� ,�  �� $�  �� $�           ,  �{ $�  �{ ,�  �� ,�  �� $�  �{ $�           ,  �� $�  �� ,�  �  ,�  �  $�  �� $�           ,  �x 0�  �x 8�  �H 8�  �H 0�  �x 0�           ,  �x @  �x !  �H !  �H @  �x @           , C @ C 8� 
� 8� 
� @ C @           ,  �  $�  �  ,� [ ,� [ $�  �  $�           , � $� � ,� @ ,� @ $� � $�           , @ $� @ ,� 8� ,� 8� $� @ $�           , (3 0� (3 8� )� 8� )� 0� (3 0�           , (3 @ (3 ! )� ! )� @ (3 @           ,      �8      �  @  �  @  �8      �8           ,  �  ��  �  ��  �  ��  �  ��  �  ��           ,  �  ��  �  �P  �  �P  �  ��  �  ��           ,  @  �8  @  �  >�  �  >�  �8  @  �8           ,  (m  ��  (m  ��  5S  ��  5S  ��  (m  ��           ,  (m  ��  (m  �P  5S  �P  5S  ��  (m  ��           ,  E�  ��  E�  ��  V�  ��  V�  ��  E�  ��           ,  >�  �8  >�  �  A�  �  A�  �8  >�  �8           ,  Z�  �8  Z�  �  ]�  �  ]�  �8  Z�  �8           ,  ]�  �8  ]�  �  }   �  }   �8  ]�  �8           ,  c�  ��  c�  ��  v�  ��  v�  ��  c�  ��           ,  c�  ��  c�  �P  v�  �P  v�  ��  c�  ��           ,  }   �8  }   �  �@  �  �@  �8  }   �8           ,  �  ��  �  ��  �>  ��  �>  ��  �  ��           ,  �  ��  �  �P  �>  �P  �>  ��  �  ��           ,      �     �  @ �  @  �      �           ,  � �  � @  � @  � �  � �           ,  �  �   �  ��  �  ��  �  �   �  �            ,  (m  �   (m @  5S @  5S  �   (m  �            ,  @  �  @ �  $� �  $�  �  @  �           ,  9;  �  9; �  >� �  >�  �  9;  �           ,  E�  �   E� @  V� @  V�  �   E�  �            ,  >�  �  >� �  A� �  A�  �  >�  �           ,  Z�  �  Z� �  ]� �  ]�  �  Z�  �           ,  c�  �   c� @  v� @  v�  �   c�  �            ,  ]�  �  ]� �  _� �  _�  �  ]�  �           ,  z�  �  z� �  }  �  }   �  z�  �           ,  �  �   � @  �> @  �>  �   �  �            ,  }   �  }  �   �    �  }   �           ,  �&  �  �& �  �@ �  �@  �  �&  �           ,  �  �@  �  ��  �  ��  �  �@  �  �@           ,      ��      �  �  �  �  ��      ��           ,  p  ��  p  �  @  �  @  ��  p  ��           ,  @  ��  @  �  >�  �  >�  ��  @  ��           ,  (m  ��  (m  ��  5S  ��  5S  ��  (m  ��           ,  (m  �@  (m  �#  5S  �#  5S  �@  (m  �@           ,  >�  ��  >�  �  ]�  �  ]�  ��  >�  ��           ,  E�  ��  E�  ��  V�  ��  V�  ��  E�  ��           ,  E�  �@  E�  �#  V�  �#  V�  �@  E�  �@           ,  c�  �@  c�  ��  v�  ��  v�  �@  c�  �@           ,  ]�  ��  ]�  �  _�  �  _�  ��  ]�  ��           ,  z�  ��  z�  �  }   �  }   ��  z�  ��           ,  �  �@  �  ��  �>  ��  �>  �@  �  �@           ,  }   ��  }   �    �    ��  }   ��           ,  �&  ��  �&  �  �@  �  �@  ��  �&  ��           ,     $�     ,�  @ ,�  @ $�     $�           ,  � 0�  � 8�  � 8�  � 0�  � 0�           ,  � @  � !  � !  � @  � @           ,  (m @  (m 8�  5S 8�  5S @  (m @           ,  @ $�  @ ,�  $� ,�  $� $�  @ $�           ,  9; $�  9; ,�  >� ,�  >� $�  9; $�           ,  E� @  E� 8�  V� 8�  V� @  E� @           ,  >� $�  >� ,�  A� ,�  A� $�  >� $�           ,  Z� $�  Z� ,�  ]� ,�  ]� $�  Z� $�           ,  c� @  c� 8�  v� 8�  v� @  c� @           ,  ]� $�  ]� ,�  _� ,�  _� $�  ]� $�           ,  z� $�  z� ,�  }  ,�  }  $�  z� $�           ,  }  $�  }  ,�  �@ ,�  �@ $�  }  $�           ,  � 0�  � 8�  �> 8�  �> 0�  � 0�           ,  � @  � !  �> !  �> @  � @           ,  �  ��  �  �   �  �   �  ��  �  ��           ,      �e      �[  �  �[  �  �e      �e           ,  p  �e  p  �[  @  �[  @  �e  p  �e           ,  @  �e  @  �[  >�  �[  >�  �e  @  �e           ,  (m  �C  (m  �   5S  �   5S  �C  (m  �C           ,  (m  ��  (m  �}  5S  �}  5S  ��  (m  ��           ,  E�  ��  E�  �   V�  �   V�  ��  E�  ��           ,  >�  �e  >�  �[  A�  �[  A�  �e  >�  �e           ,  Z�  �e  Z�  �[  ]�  �[  ]�  �e  Z�  �e           ,  ]�  �e  ]�  �[  }   �[  }   �e  ]�  �e           ,  c�  �C  c�  �   v�  �   v�  �C  c�  �C           ,  c�  ��  c�  �}  v�  �}  v�  ��  c�  ��           ,  �  ��  �  �   �>  �   �>  ��  �  ��           ,  }   �e  }   �[    �[    �e  }   �e           ,  �&  �e  �&  �[  �@  �[  �@  �e  �&  �e           ,  �      �  @  �  @  �      �               ,      �      �  �  �  �  �      �           ,  p  �  p  �  @  �  @  �  p  �           ,  @  �  @  �  >�  �  >�  �  @  �           ,  (m  p  (m  @  5S  @  5S  p  (m  p           ,  (m      (m  �  5S  �  5S      (m               ,  >�  �  >�  �  ]�  �  ]�  �  >�  �           ,  E�  p  E�  @  V�  @  V�  p  E�  p           ,  E�      E�  �  V�  �  V�      E�               ,  ]�  �  ]�  �  }   �  }   �  ]�  �           ,  c�  p  c�  @  v�  @  v�  p  c�  p           ,  c�      c�  �  v�  �  v�      c�               ,  }   �  }   �  �@  �  �@  �  }   �           ,  �  p  �  @  �>  @  �>  p  �  p           ,  �      �  �  �>  �  �>      �               ,      %�      7�  @  7�  @  %�      %�           ,  �  ;�  �  >�  �  >�  �  ;�  �  ;�           ,  �  @  �  !�  �  !�  �  @  �  @           ,  (m  @  (m  >�  5S  >�  5S  @  (m  @           ,  @  %�  @  7�  $�  7�  $�  %�  @  %�           ,  9;  %�  9;  7�  >�  7�  >�  %�  9;  %�           ,  E�  @  E�  >�  V�  >�  V�  @  E�  @           ,  >�  %�  >�  7�  A�  7�  A�  %�  >�  %�           ,  Z�  %�  Z�  7�  ]�  7�  ]�  %�  Z�  %�           ,  ]�  %�  ]�  7�  }   7�  }   %�  ]�  %�           ,  c�  ;�  c�  >�  v�  >�  v�  ;�  c�  ;�           ,  c�  @  c�  !�  v�  !�  v�  @  c�  @           ,  }   %�  }   7�  �@  7�  �@  %�  }   %�           ,  �  ;�  �  >�  �>  >�  �>  ;�  �  ;�           ,  �  @  �  !�  �>  !�  �>  @  �  @           ,  �  >�  �  ]�  �  ]�  �  >�  �  >�           ,      E%      W  �  W  �  E%      E%           ,  p  E%  p  W  @  W  @  E%  p  E%           ,  @  E%  @  W  >�  W  >�  E%  @  E%           ,  (m  [  (m  ]�  5S  ]�  5S  [  (m  [           ,  (m  >�  (m  A=  5S  A=  5S  >�  (m  >�           ,  E�  >�  E�  ]�  V�  ]�  V�  >�  E�  >�           ,  >�  E%  >�  W  A�  W  A�  E%  >�  E%           ,  Z�  E%  Z�  W  ]�  W  ]�  E%  Z�  E%           ,  ]�  E%  ]�  W  }   W  }   E%  ]�  E%           ,  c�  [  c�  ]�  v�  ]�  v�  [  c�  [           ,  c�  >�  c�  A=  v�  A=  v�  >�  c�  >�           ,  �  >�  �  ]�  �>  ]�  �>  >�  �  >�           ,  }   E%  }   W    W    E%  }   E%           ,  �&  E%  �&  W  �@  W  �@  E%  �&  E%           ,      ix      qH  @  qH  @  ix      ix           ,  �  u0  �  }   �  }   �  u0  �  u0           ,  �  ]�  �  e�  �  e�  �  ]�  �  ]�           ,  @  ix  @  qH  >�  qH  >�  ix  @  ix           ,  (m  u0  (m  }   5S  }   5S  u0  (m  u0           ,  (m  ]�  (m  e�  5S  e�  5S  ]�  (m  ]�           ,  E�  ]�  E�  }   V�  }   V�  ]�  E�  ]�           ,  >�  ix  >�  qH  A�  qH  A�  ix  >�  ix           ,  Z�  ix  Z�  qH  ]�  qH  ]�  ix  Z�  ix           ,  c�  ]�  c�  }   v�  }   v�  ]�  c�  ]�           ,  ]�  ix  ]�  qH  _�  qH  _�  ix  ]�  ix           ,  z�  ix  z�  qH  }   qH  }   ix  z�  ix           ,  �  ]�  �  }   �>  }   �>  ]�  �  ]�           ,  }   ix  }   qH    qH    ix  }   ix           ,  �&  ix  �&  qH  �@  qH  �@  ix  �&  ix           ,      �u      ��  @  ��  @  �u      �u           ,  �  �]  �  �@  �  �@  �  �]  �  �]           ,  �  }   �  ��  �  ��  �  }   �  }            ,  @  �u  @  ��  >�  ��  >�  �u  @  �u           ,  (m  �]  (m  �@  5S  �@  5S  �]  (m  �]           ,  (m  }   (m  ��  5S  ��  5S  }   (m  }            ,  E�  }   E�  �@  V�  �@  V�  }   E�  }            ,  >�  �u  >�  ��  A�  ��  A�  �u  >�  �u           ,  Z�  �u  Z�  ��  ]�  ��  ]�  �u  Z�  �u           ,  ]�  �u  ]�  ��  }   ��  }   �u  ]�  �u           ,  c�  �]  c�  �@  v�  �@  v�  �]  c�  �]           ,  c�  }   c�  ��  v�  ��  v�  }   c�  }            ,  }   �u  }   ��  �@  ��  �@  �u  }   �u           ,  �  �]  �  �@  �>  �@  �>  �]  �  �]           ,  �  }   �  ��  �>  ��  �>  }   �  }            ,  �@  E%  �@  W  ��  W  ��  E%  �@  E%           ,  �c  [  �c  ]�  �]  ]�  �]  [  �c  [           ,  �c  >�  �c  A=  �]  A=  �]  >�  �c  >�           ,  ��  E%  ��  W  ��  W  ��  E%  ��  E%           ,  ĭ  [  ĭ  ]�  ѓ  ]�  ѓ  [  ĭ  [           ,  ĭ  >�  ĭ  A=  ѓ  A=  ѓ  >�  ĭ  >�           ,  �x  >�  �x  ]�  �H  ]�  �H  >�  �x  >�           ,  ��  E%  ��  W  �  W  �  E%  ��  E%           ,  �0  E%  �0  W  �   W  �   E%  �0  E%           ,  �   E%  �   W @  W @  E%  �   E%           , C  [ C  ]� 
�  ]� 
�  [ C  [           , C  >� C  A= 
�  A= 
�  >� C  >�           , @  E% @  W 8�  W 8�  E% @  E%           , (3  [ (3  ]� )�  ]� )�  [ (3  [           , (3  >� (3  A= )�  A= )�  >� (3  >�           ,  �@  %�  �@  7�  ��  7�  ��  %�  �@  %�           ,  �c  ;�  �c  >�  �]  >�  �]  ;�  �c  ;�           ,  �c  @  �c  !�  �]  !�  �]  @  �c  @           ,  ĭ  @  ĭ  >�  ѓ  >�  ѓ  @  ĭ  @           ,  ��  %�  ��  7�  ��  7�  ��  %�  ��  %�           ,  �{  %�  �{  7�  ��  7�  ��  %�  �{  %�           ,  �x  @  �x  >�  �H  >�  �H  @  �x  @           ,  ��  %�  ��  7�  �  7�  �  %�  ��  %�           ,  �0  %�  �0  7�  �   7�  �   %�  �0  %�           ,  �   %�  �   7� @  7� @  %�  �   %�           , C  ;� C  >� 
�  >� 
�  ;� C  ;�           , C  @ C  !� 
�  !� 
�  @ C  @           , @  %� @  7� 8�  7� 8�  %� @  %�           , (3  ;� (3  >� )�  >� )�  ;� (3  ;�           , (3  @ (3  !� )�  !� )�  @ (3  @           ,  �c  ]�  �c  }   �]  }   �]  ]�  �c  ]�           ,  �@  ix  �@  qH  �{  qH  �{  ix  �@  ix           ,  �E  ix  �E  qH  ��  qH  ��  ix  �E  ix           ,  ��  ix  ��  qH  ��  qH  ��  ix  ��  ix           ,  ĭ  u0  ĭ  }   ѓ  }   ѓ  u0  ĭ  u0           ,  ĭ  ]�  ĭ  e�  ѓ  e�  ѓ  ]�  ĭ  ]�           ,  ��  ix  ��  qH  �   qH  �   ix  ��  ix           ,  �x  u0  �x  }   �H  }   �H  u0  �x  u0           ,  �x  ]�  �x  e�  �H  e�  �H  ]�  �x  ]�           , C  ]� C  }  
�  }  
�  ]� C  ]�           ,  �   ix  �   qH [  qH [  ix  �   ix           , �  ix �  qH @  qH @  ix �  ix           , @  ix @  qH 8�  qH 8�  ix @  ix           , (3  u0 (3  }  )�  }  )�  u0 (3  u0           , (3  ]� (3  e� )�  e� )�  ]� (3  ]�           ,  �@  �  �@  �  ��  �  ��  �  �@  �           ,  �c  p  �c  @  �]  @  �]  p  �c  p           ,  �c      �c  �  �]  �  �]      �c               ,  ĭ      ĭ  @  ѓ  @  ѓ      ĭ               ,  ��  �  ��  �  ��  �  ��  �  ��  �           ,  �{  �  �{  �  ��  �  ��  �  �{  �           ,  ��  �  ��  �  �   �  �   �  ��  �           ,  �x  p  �x  @  �H  @  �H  p  �x  p           ,  �x      �x  �  �H  �  �H      �x               ,  �   �  �   � @  � @  �  �   �           , C  p C  @ 
�  @ 
�  p C  p           , C     C  � 
�  � 
�     C               , (3     (3  @ )�  @ )�     (3               , @  � @  � %�  � %�  � @  �           , ,  � ,  � 8�  � 8�  � ,  �           ,  �c  }   �c  �@  �]  �@  �]  }   �c  }            ,  �@  �u  �@  ��  �{  ��  �{  �u  �@  �u           ,  �E  �u  �E  ��  ��  ��  ��  �u  �E  �u           ,  ��  �u  ��  ��  ��  ��  ��  �u  ��  �u           ,  ĭ  �]  ĭ  �@  ѓ  �@  ѓ  �]  ĭ  �]           ,  ĭ  }   ĭ  ��  ѓ  ��  ѓ  }   ĭ  }            ,  ��  �u  ��  ��  �   ��  �   �u  ��  �u           ,  �x  �]  �x  �@  �H  �@  �H  �]  �x  �]           ,  �x  }   �x  ��  �H  ��  �H  }   �x  }            , C  }  C  �@ 
�  �@ 
�  }  C  }            ,  �   �u  �   �� [  �� [  �u  �   �u           , �  �u �  �� @  �� @  �u �  �u           , (3  }  (3  �@ )�  �@ )�  }  (3  }            , @  �u @  �� %�  �� %�  �u @  �u           , ,  �u ,  �� 8�  �� 8�  �u ,  �u      