VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO my_logo
  CLASS BLOCK ;
  FOREIGN my_logo ;
  SIZE 32.000 BY 32.000 ;
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 0.000 8.000 1.500 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 24.000 0.000 32.000 1.500 ;
    END
  END VGND
  OBS
      LAYER Metal1 ;
        RECT 0.000 4.000 32.000 32.000 ;
      LAYER Metal2 ;
        RECT 0.000 4.000 32.000 32.000 ;
      LAYER Metal3 ;
        RECT 0.000 4.000 32.000 32.000 ;
      LAYER Metal4 ;
        RECT 0.000 4.000 32.000 32.000 ;
  END
END my_logo
END LIBRARY
