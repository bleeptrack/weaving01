# LEF file generated for my_logo
VERSION 5.8 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO my_logo
   CLASS BLOCK ;
   FOREIGN my_logo 0 0 ;
   SIZE 32.000 BY 32.000 ;
   SYMMETRY X Y ;
   PIN VDD
      DIRECTION INOUT ;
      USE POWER ;
      PORT
         LAYER Metal1 ;
         RECT 0.000 30.000 32.000 32.000 ;
      END
   END VDD
   PIN VSS
      DIRECTION INOUT ;
      USE GROUND ;
      PORT
         LAYER Metal1 ;
         RECT 0.000 0.000 32.000 2.000 ;
      END
   END VSS
   PIN in
      DIRECTION INPUT ;
      USE SIGNAL ;
      PORT
         LAYER Metal1 ;
         RECT 0.000 14.000 2.000 18.000 ;
      END
   END in
   PIN out
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      PORT
         LAYER Metal1 ;
         RECT 30.000 14.000 32.000 18.000 ;
      END
   END out
   OBS
      LAYER Metal1 ;
      RECT 0.000 0.000 32.000 32.000 ;
   END
END my_logo
