# LEF file generated for my_logo
VERSION 5.8 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO my_logo
   CLASS BLOCK ;
   FOREIGN my_logo 0 0 ;
   SIZE 80.000 BY 80.000 ;
   SYMMETRY X Y ;
   OBS
      LAYER Metal1 ;
      RECT 0.000 0.000 80.000 80.000 ;
   END
END my_logo
